# Input constraints
set_property PACKAGE_PIN AA12 [get_ports {a[0]}]
set_property PACKAGE_PIN AA13 [get_ports {a[1]}]
set_property PACKAGE_PIN AA14 [get_ports {a[2]}]
set_property PACKAGE_PIN AA15 [get_ports {a[3]}]

set_property PACKAGE_PIN AB12 [get_ports {b[0]}]
set_property PACKAGE_PIN AB13 [get_ports {b[1]}]
set_property PACKAGE_PIN AB14 [get_ports {b[2]}]
set_property PACKAGE_PIN AB15 [get_ports {b[3]}]

set_property PACKAGE_PIN AC12 [get_ports c_in]

# Output constraints
set_property PACKAGE_PIN AD12 [get_ports {sum[0]}]
set_property PACKAGE_PIN AD13 [get_ports {sum[1]}]
set_property PACKAGE_PIN AD14 [get_ports {sum[2]}]
set_property PACKAGE_PIN AD15 [get_ports {sum[3]}]

set_property PACKAGE_PIN AE12 [get_ports GG]
set_property PACKAGE_PIN AE13 [get_ports GP]
set_property PACKAGE_PIN AE14 [get_ports c_out]
